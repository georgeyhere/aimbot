module cam_capture_maxis_tb();


endmodule
